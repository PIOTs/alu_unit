----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    12:16:13 09/25/2015 
-- Design Name: 
-- Module Name:    arithm_unit - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity arithm_unit is
port(i_a:in std_logic_vector(31 downto 0);
	  i_b:in std_logic_vector(31 downto 0);
	  cin:in std_logic;
	  s:in std_logic_vector(1 downto 0);
	  result:out std_logic_vector(32 downto 0));
end arithm_unit;

architecture Behavioral of arithm_unit is

	component mux_4to1 is
	port(a,b,c,d:in std_logic;
		s:in std_logic_vector(1 downto 0);
		y:out std_logic);
	end component;
	
	component addr_32bit is
	port(i_a:in std_logic_vector(31 downto 0);
	  i_b:in std_logic_vector(31 downto 0);
	  cin:in std_logic;
	  result:out std_logic_vector(32 downto 0));
	end component;
  
  signal sg:std_logic_vector(31 downto 0);----signal generated by 4:1_1bit mux e.g Y0,Y1,Y2...etc  

begin

p0:mux_4to1 port map(i_b(0),not i_b(0),'1','0',s,sg(0));
p1:mux_4to1 port map(i_b(1),not i_b(1),'1','0',s,sg(1));
p2:mux_4to1 port map(i_b(2),not i_b(2),'1','0',s,sg(2));
p3:mux_4to1 port map(i_b(3),not i_b(3),'1','0',s,sg(3));
p4:mux_4to1 port map(i_b(4),not i_b(4),'1','0',s,sg(4));
p5:mux_4to1 port map(i_b(5),not i_b(5),'1','0',s,sg(5));
p6:mux_4to1 port map(i_b(6),not i_b(6),'1','0',s,sg(6));
p7:mux_4to1 port map(i_b(7),not i_b(7),'1','0',s,sg(7));
p8:mux_4to1 port map(i_b(8),not i_b(8),'1','0',s,sg(8));
p9:mux_4to1 port map(i_b(9),not i_b(9),'1','0',s,sg(9));
p10:mux_4to1 port map(i_b(10),not i_b(10),'1','0',s,sg(10));
p11:mux_4to1 port map(i_b(11),not i_b(11),'1','0',s,sg(11));
p12:mux_4to1 port map(i_b(12),not i_b(12),'1','0',s,sg(12));
p13:mux_4to1 port map(i_b(13),not i_b(13),'1','0',s,sg(13));
p14:mux_4to1 port map(i_b(14),not i_b(14),'1','0',s,sg(14));
p15:mux_4to1 port map(i_b(15),not i_b(15),'1','0',s,sg(15));
p16:mux_4to1 port map(i_b(16),not i_b(16),'1','0',s,sg(16));
p17:mux_4to1 port map(i_b(17),not i_b(17),'1','0',s,sg(17));
p18:mux_4to1 port map(i_b(18),not i_b(18),'1','0',s,sg(18));
p19:mux_4to1 port map(i_b(19),not i_b(19),'1','0',s,sg(19));
p20:mux_4to1 port map(i_b(20),not i_b(20),'1','0',s,sg(20));
p21:mux_4to1 port map(i_b(21),not i_b(21),'1','0',s,sg(21));
p22:mux_4to1 port map(i_b(22),not i_b(22),'1','0',s,sg(22));
p23:mux_4to1 port map(i_b(23),not i_b(23),'1','0',s,sg(23));
p24:mux_4to1 port map(i_b(24),not i_b(24),'1','0',s,sg(24));
p25:mux_4to1 port map(i_b(25),not i_b(25),'1','0',s,sg(25));
p26:mux_4to1 port map(i_b(26),not i_b(26),'1','0',s,sg(26));
p27:mux_4to1 port map(i_b(27),not i_b(27),'1','0',s,sg(27));
p28:mux_4to1 port map(i_b(28),not i_b(28),'1','0',s,sg(28));
p29:mux_4to1 port map(i_b(29),not i_b(29),'1','0',s,sg(29));
p30:mux_4to1 port map(i_b(30),not i_b(30),'1','0',s,sg(30));
p31:mux_4to1 port map(i_b(31),not i_b(31),'1','0',s,sg(31));

p32:addr_32bit port map(i_a,sg,cin,result);


end Behavioral;

